***6T SRAM READ MODE***

.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7

.subckt inverter in out vdd
M1 out in vdd vdd pmod w=100u l=10u
M2 out in 0 0 nmod w=100u l=10u
.ends inverter

Vdd 2 0 dc 5

Vwl 6 0 dc 5

.IC V(3)=5

Xq 3 1 2 inverter
Xqbar 1 3 2 inverter

M5 7 6 3 3 nmod w=100u l=10u
M6 8 6 1 1 nmod w=100u l=10u

C7 7 0 1u IC=2.5
C8 8 0 1u IC=2.5

.tran 0.1m 400m
.control
run
plot v(7) v(8) v(3) v(1)
.endc
.end